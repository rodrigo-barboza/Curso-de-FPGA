LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DISP_CONTROL IS PORT (
	BAR: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
	CLK:  IN STD_LOGIC
);
END DISP_CONTROL;

ARCHITECTURE DISP_CONTROL_HW OF DISP_CONTROL IS BEGIN
	PROCESS (CLK) 
		-- VARIÁVEL PARA CONTAR DE 0 ATÉ 10, DO TIPO INTEIRO
		-- VARIÁVEL DE NOME "COUNTER" DO TIPO INTEIRO E QUE CONTA DE 0 ATÉ 10
		VARIABLE COUNTER: INTEGER RANGE 0 TO 10;
	BEGIN
		IF (CLK = '1') THEN
			-- ATRIBUIÇÃO DE VARIÁVEIS É FEITA COM := E NÃO COM <=
			COUNTER := COUNTER + 1;
			
			IF (COUNTER = 10) THEN
				COUNTER := 0;
			END IF;
		END IF;
		
		CASE COUNTER IS 
			WHEN 0 => BAR <= "1111110";
			WHEN 1 => BAR <= "0110000";
			WHEN 2 => BAR <= "1100111";
			WHEN 3 => BAR <= "0001110";
			WHEN 4 => BAR <= "0011010";
			WHEN 5 => BAR <= "1101010";
			WHEN 6 => BAR <= "0110101";
			WHEN 7 => BAR <= "1010101";
			WHEN 8 => BAR <= "0101010";
			WHEN 9 => BAR <= "1001100";
			WHEN OTHERS => BAR <= "0000000";
		END CASE;
	END PROCESS;
END DISP_CONTROL_HW;
	