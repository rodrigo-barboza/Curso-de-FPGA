ENTITY TESTBENCH1 IS END; -- O TB1 � UMA ENTIDADE SEM ENTRADAS OU SA�DAS.

-- BIBLI�TECAS E PACOTES
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE STD.TEXTIO.ALL;

ARCHITECTURE XOR_GATE_TB OF TESTBENCH1 IS 
COMPONENT XOR_GATE PORT (
  A:  IN STD_LOGIC;
  B:  IN STD_LOGIC;
  C: OUT STD_LOGIC
); 
END COMPONENT;
  -- SINAIS AUXILIARES PARA INTERCONEX�O AO PROCESSO DE ESTIMULO
  SIGNAL I_1: STD_LOGIC;
  SIGNAL I_2: STD_LOGIC;
  -- C�DIGO CONCORRENTE
BEGIN
  -- CRIAR INST�NCIA DO COMPONENTE XOR_GATE PARA INTERCONEX�O DO COMPONENTE COM O PROCESSO DE ESTIMULO
  XOR1: XOR_GATE PORT MAP (A => I_1, B => I_2, C => OPEN);
    ESTIMULO: PROCESS BEGIN
      WAIT FOR 5 NS; I_1 <= '0'; I_2 <= '0';
      WAIT FOR 5 NS; I_1 <= '1';
      WAIT FOR 5 NS; I_2 <= '1';
      WAIT FOR 5 NS; I_1 <= '0';
      WAIT;
    END PROCESS ESTIMULO;
END XOR_GATE_TB;
      