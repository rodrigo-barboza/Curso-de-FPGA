-- AUTOR: RODRIGO BARBOZA
-- DATA: 31/03/2020

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY XOR_GATE IS PORT (
  A: IN  STD_LOGIC;
  B: IN  STD_LOGIC;
  C: OUT STD_LOGIC
);
END XOR_GATE;

ARCHITECTURE XOR_GATE_HW OF XOR_GATE IS BEGIN
  C <= A XOR B;
END XOR_GATE_HW;
