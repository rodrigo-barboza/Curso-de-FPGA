LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX_4b IS PORT (
	SEL: IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
	  A: IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
	  X: OUT STD_LOGIC
);
END MUX_4b;

ARCHITECTURE MUX_4b_HARD OF MUX_4b IS
BEGIN
	WITH SEL SELECT
		X <= A(0) WHEN "00",
			  A(1) WHEN "10",
			  A(2) WHEN "01",
			  A(3) WHEN "11",
			  '0' when others;
	
END MUX_4b_HARD;
